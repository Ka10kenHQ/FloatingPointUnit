module muldiv (
    input sa,
    input sb,
    input [52:0] fa,
    input [52:0] fb,
    input [10:0] ea,
    input [10:0] eb,
    input [5:0] lza,
    input [5:0] lzb,
    input [52:0] nan,
    input [3:0] fla,
    input [3:0] flb,
    output reg [56:0] fq,
    output reg [12:0] eq,
    output reg sq,
    output reg [3:0] flq
);


endmodule
