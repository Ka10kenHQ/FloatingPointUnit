module tb_ftadd;

  parameter n = 13;
  
  reg [n-1:0] a;
  reg [n-1:0] b;
  reg [n-1:0] c;
  reg [n-1:0] d;

  wire [n:0] t;
  wire [n:0] s;

  ftadd #(n) uut (
      .a(a),
      .b(b),
      .c(c),
      .d(d),
      .t(t),
      .s(s)
  );

  initial begin
    $monitor("Time = %0t | a = %d, b = %d, c = %d, d = %d | t = %d, s = %d", $time, a, b, c, d, t, s);

    a = 13'b0000000000001; 
    b = 13'b0000000000010; 
    c = 13'b0000000000100;
    d = 13'b0000000001000;

    #10 a = 13'b0101010101010; b = 13'b1100110011001; c = 13'b1010101010101; d = 13'b0011001100110;
    #10 a = 13'b1111111111111; b = 13'b0000000000000; c = 13'b0000000001111; d = 13'b1010101010101;
    #10 a = 13'b1001100110011; b = 13'b0101010101010; c = 13'b1110000000000; d = 13'b0001111100000;
    #10 a = 13'b0001110001110; b = 13'b1111111111111; c = 13'b0000000000000; d = 13'b1111000001110;
    #10 a = 13'b1101010101010; b = 13'b1110000001110; c = 13'b1010101010101; d = 13'b0000000000001;

  end

endmodule

