module normshift(
    input [56:0] fr,
    input [12:0] er,
    input OVFen,
    input UNFen,

    output [127:0] fn,
    output [10:0] eni,
    output [10:0] en,
    output TINY,
    output OVF1
);




endmodule
