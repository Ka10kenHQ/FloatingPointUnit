module multree(
    input [57:0] a,
    input [57:0] b,

    output [115:0] out
);


endmodule
