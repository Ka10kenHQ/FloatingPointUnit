module inf_selector (
    input [1:0] RM,
    input s,
    output inf
);


endmodule

