module tb_unpacker;

    parameter N = 64;
    
    reg dbs;
    reg [N-1:0] x;
    reg ez;
    reg normal;

    wire [5:0] lz;
    wire [52:0] f;
    wire fz;
    wire [51:0] h;

    unpacker #(N) uut (
        .dbs(dbs),
        .x(x),
        .ez(ez),
        .normal(normal),
        .lz(lz),
        .f(f),
        .fz(fz),
        .h(h)
    );

    initial begin
        dbs = 0;
        x = 64'hA5A5A5A5A5A5A5A5;  // Sample input value
        ez = 0;
        normal = 1;
        #10;
        
        dbs = 1;
        x = 64'h1F1F1F1F1F1F1F1F;  // Another sample input value
        ez = 1;
        normal = 0;
        #10;

        dbs = 0;
        x = 64'hDEADBEEFDEADBEEF;  // Another input pattern
        ez = 0;
        normal = 1;
        #10;

        dbs = 1;
        x = 64'hFFFFFFFFFFFFFFFF;  // All bits set
        ez = 1;
        normal = 0;
        #10;

        dbs = 0;
        x = 64'h1234567890ABCDEF;  // Random 64-bit value
        ez = 0;
        normal = 1;
        #10;

        $finish;  
    end

    initial begin
        $monitor("At time %t, dbs = %b, x = %h, ez = %b, normal = %b, lz = %h, f = %h, fz = %b, h = %h", 
                  $time, dbs, x, ez, normal, lz, f, fz, h);
    end

endmodule
