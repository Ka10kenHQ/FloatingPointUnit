module exprnd(
    input s,
    input [10:0] e3,
    input [52:0] f3,
    input [1:0] RM,
    input OVF,
    input db,
    input OVFen,

    output [10:0] eout,
    output [51:0] fout
);

wire inf;
assign inf = (RM[1] == 1'b1) ? RM[0] : ~(RM[0] ^ s);

assign eout = (OVF & ~OVFen) ? 
              (inf ? {{3{db}}, 8'b11111111} : {{3{db}}, 7'b1111111, 1'b0}) :
              (e3 & f3[52]);

assign fout = (OVF & ~OVFen) ? 
              (inf ? 52'b0 : {{23{1'b1}}, {29{db}}}) :
              f3[51:0];

endmodule

