module div_logic(
    input           clk,
    input           rst_n,
    input  [52:0]   fa,
    input  [52:0]   fb,
    input           db,
    input           fdiv,
    output logic [56:0] fq
);

logic  [57:0] fa_in, fb_in;
logic [115:0] mul_out;
wire [56:0] fd_out;
logic or_out;
logic [7:0] rom_data;
parameter n = 60;

logic [3:0] state;
logic [1:0] Dcnt;
logic [57:0] x, A, Da, Db;
logic [54:0] E;
logic [115:0] Eb;
logic [8:0] look_up;

rom256X8 rom_inst (.addr(fb[51:44]), .data(rom_data));
multree mlt (.a(fa_in), .b(fb_in), .out(mul_out));
ortree #(n) or_inst (.x(mul_out[59:0]), .or_out(or_out));
select_fd_reg fd_inst_reg (
    .clk(clk),
    .Da(Da),
    .Db(Db),
    .Eb(Eb[114:0]),
    .E(E),
    .db(db),
    .fd(fd_out)
);

localparam IDLE    = 4'd0;
localparam NEWTON1 = 4'd1;
localparam NEWTON2 = 4'd2;
localparam NEWTON3 = 4'd3;
localparam NEWTON4 = 4'd4;
localparam QUOT1   = 4'd5;
localparam QUOT2   = 4'd6;
localparam QUOT3   = 4'd7;
localparam QUOT4   = 4'd8;
localparam RESULT  = 4'd9;

always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        state <= IDLE;
        Dcnt  <= 0;
        x     <= 0;
        A     <= 0;
        Da    <= 0;
        Db    <= 0;
        E     <= 0;
        Eb    <= 0;
        fa_in <= 0;
        fb_in <= 0;
        fq    <= 0;
        look_up <= 0;
    end else begin
        case (state)
            IDLE: begin
                look_up <= rom_data;
                x       <= {2'b01, rom_data, 48'b0};
                Dcnt    <= db ? 2'b11 : 2'b10;
                state   <= NEWTON1;
            end

            NEWTON1: begin
                fa_in <= x;
                fb_in <= {fb[51:0], 6'b0};
                Dcnt  <= Dcnt - 1;
                state <= NEWTON2;
            end

            NEWTON2: begin
                A     <= ~mul_out[115:58];
                state <= NEWTON3;
            end

            NEWTON3: begin
                fa_in <= A;
                fb_in <= x;
                state <= NEWTON4;
            end

            NEWTON4: begin
                x <= mul_out[115:58];
                if (Dcnt == 2'b00)
                    state <= QUOT1;
                else
                    state <= NEWTON1;
            end

            QUOT1: begin
                fa_in <= {fa[51:0], 6'b0};
                fb_in <= x;
                state <= QUOT2;
            end

            QUOT2: begin
                Da <= {fa,5'b0};
                Db <= {fb,5'b0};
                E  <= {mul_out[115:90], mul_out[89:61] & {29{db}}};
                Eb <= mul_out;
                state <= QUOT3;
            end

            QUOT3: begin
                state <= RESULT;
            end

            RESULT: begin
                fq <= fd_out;
                state <= RESULT;
            end
        endcase
    end
end

endmodule
