module sigfmd (
    input [52:0] fa,
    input [52:0] fb,
    output reg [56:0] fq
);



endmodule
