Module RoundingModes #(parameter NUM_REGS = 4, 
parameter DEPTH = 4 // Number of rounding modes
) (


);

logic [WIDTH-1:0] reg_file [0:]




endmodule