module adder(
    input [52:0] fa,
    input [10:0] ea,
    input sa,
    input [52:0] fb,
    input [10:0] eb,
    input sb,
    input sub,
    input fla,
    input flb,
    input nan
    );

endmodule
