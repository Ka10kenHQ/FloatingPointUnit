module sigfmd (
    input [52:0] fa,
    input [52:0] fb,
    input fdiv,
    input tlu,
    input db,
    output reg [56:0] fq
);




endmodule
