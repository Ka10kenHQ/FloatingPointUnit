module master  (
);


// TODO

endmodule
