module expnorm(
    input [10:0] er,
    input [5:0] lz,

    input db,
    input OVFen,
    input OVF1,
    input UNFen,
    input TINY,


    output [10:0] eni,
    output [10:0] en
);


endmodule
