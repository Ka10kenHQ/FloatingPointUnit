module alignment(
    input [10:0] ea,
    input [10:0] eb,

    input [52:0] fa,
    input  sa,
    
    input [52:0] fb,
    input  sb,
    
    output reg[10:0] es,
    output reg[55:0] fb3,
    output [52:0] fa2,
    output  sa2,
    output reg sx,
    output  sb2
);

wire [10:0] as;
wire eb_gt_ea;

exp_sub uut(
    .ea(ea),
    .eb(eb),
    .as(as),
    .eb_gt_ea(eb_gt_ea)
);

wire [5:0] as2;

limit uut1(
    .as(as),
    .eb_gt_ea(eb_gt_ea),
    .as2(as2)
);

wire [54:0] fb2;
swap uut2(
    .fa(fa),
    .fb(fb),
    .sa(sa),
    .sb(sb),
    .eb_gt_ea(eb_gt_ea),
    .fb2(fb2),
    .fa2(fa2),
    .sa2(sa2),
    .sb2(sb2)
);

wire [54:0] fp3_h;

lrs uut3(
.as2(as2),
.fb2(fb2),
.fb3(fp3_h)
);

wire sticky;
sticky uut4(
.as2(as2),
.fb2(fb2),
.sticky(sticky)
);

always@(*) begin
sx = sa2 ^ sb2;
es = eb_gt_ea ? eb : ea;
fb3 = {fp3_h[54:0], sticky};
end    
endmodule
