module master  (
);

// TODO

endmodule
