module signormshift(
    input [56:0] fr,
    input [12:0] sh,

    output [127:0] fn
);



endmodule
