module signormshift(

);



endmodule
