module alignment (
    input [10:0] ea,
    input [10:0] eb,
    input [52:0] fa,
    input sa,
    input [52:0] fb,
    input sb
    );


endmodule
