`include "./../tb_spec"
module tb_spec;

    reg sb;
    reg sa;
    reg [52:0] fla;
    reg [52:0] flb;
    wire INFs;
    wire NANs;
    wire INV;

    spec uut (
        .sb(sb),
        .sa(sa),
        .fla(fla),
        .flb(flb),
        .INFs(INFs),
        .NANs(NANs),
        .INV(INV)
    );

    initial begin
        sb = 0; sa = 0; fla = 53'b0; flb = 53'b0;
        #10 sb = 1; sa = 1; fla = 53'b10000000000000000000000000000000000000000000000000000; flb = 53'b10000000000000000000000000000000000000000000000000000;
        #10 sb = 0; sa = 1; fla = 53'b11000000000000000000000000000000000000000000000000000; flb = 53'b00100000000000000000000000000000000000000000000000000;
        #10 sb = 1; sa = 0; fla = 53'b00010000000000000000000000000000000000000000000000000; flb = 53'b11100000000000000000000000000000000000000000000000000;
        #10 sb = 1; sa = 1; fla = 53'b00000000000000000000000000000000000000000000000000000; flb = 53'b10000000000000000000000000000000000000000000000000000;
        #10 sb = 0; sa = 0; fla = 53'b11111111111111111111111111111111111111111111111111111; flb = 53'b01111111111111111111111111111111111111111111111111111;
        #10 sb = 0; sa = 1; fla = 53'b01000000000000000000000000000000000000000000000000000; flb = 53'b00000000000000000000000000000000000000000000000000000;
        #10 sb = 1; sa = 0; fla = 53'b00100000000000000000000000000000000000000000000000000; flb = 53'b10000000000000000000000000000000000000000000000000000;
        #10;
    end

endmodule

