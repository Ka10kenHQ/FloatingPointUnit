module Master #(parameter WIDTH = 64) (
    input logic [WIDTH-1:0] FA2,
    input logic [WIDTH-1:0] FB2
);
always_comb begin
    
end

endmodule