module adder(
    input [52:0] fa,
    input [10:0] ea,
    input sa,
    input [52:0] fb,
    input [10:0] eb,
    input sb,
    input sub,
    input fla,
    input flb,
    input nan,
    output [10:0] es,
    output [56:0] fs,
    output ss,
    output fls
    );

endmodule
