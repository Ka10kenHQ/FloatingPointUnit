module tb_lrs;

    reg [6:0] as2;
    reg [54:0] fb2;
    wire [54:0] fb3;

    lrs uut (
        .as2(as2),
        .fb2(fb2),
        .fb3(fb3)
    );

    initial begin
        $display("Time | as2     | fb2                                         | fb3");
        $monitor("%4t | %b      | %b | %b", $time, as2, fb2, fb3);

        as2 = 7'b1010101; fb2 = 55'b110110101101110101101110101101110101101110110110101101110101101; #10;
        as2 = 7'b0000000; fb2 = 55'b1010101010101010101010101010101010101010101010101010101010101010; #10;
        as2 = 7'b1111111; fb2 = 55'b001100110011001100110011001100110011001100110011001100110011001; #10;
        as2 = 7'b1011101; fb2 = 55'b010101010101010101010101010101010101010101010101010101010101010; #10;
        as2 = 7'b0001101; fb2 = 55'b111111111111111111111111111111111111111111111111111111111111111; #10;
        
        $stop;
    end

endmodule

